/*=================================================================================================
 = File name : ALU_seqr.sv                                                                        =
 = Author    : Sherif Omar                                                                        =
 = Linkedin  : https://www.linkedin.com/in/sherif-omar-23829b222/                                 =
 = Email     : sherifomar661@gmail.com  "If you have any questions, feel free to contact me"      =
 = Date      : Sep 09 , 2022                                                                      =
 =================================================================================================*/

`ifndef ALU_SEQR
`define ALU_SEQR
typedef uvm_sequencer#(ALU_trans) ALU_seqr;
`endif